`timescale 1ns/100ps
`include "sort_reg.v"

`define CYCLE 10

module tb_sort_reg;
  
  reg  [4:0] old_index;
  reg  [28:0] Q;
  reg clk, reset;
  
  //wire [31:0] asi;
  wire [28:0] s1, s2, s3, s4, s5, s6, s7, s8, s9, s10, s11, s12, s13, s14, s15, s16, s17, s18, s19, s20, s21, s22, s23, s24, s25, s26, s27, s28, s29, s30, s31, s32;

sort_reg sr(old_index, Q, clk, reset, s1, s2, s3, s4, s5, s6, s7, s8, s9, s10, s11, s12, s13, s14, s15, s16,
 s17, s18, s19, s20, s21, s22, s23, s24, s25, s26, s27, s28, s29, s30, s31, s32);


//initial $sdf_annotate("sorting.sdf", sr);

  always #(`CYCLE/2) clk = ~clk;

  initial
  begin
    reset=1; clk=1;
    #5 reset=0;
    #10 old_index=5'b00000 ; Q=29'b00000_00_000001_00000010_00000010; 
    #10 old_index=5'b00001 ; Q=29'b00001_00_000001_00000010_00010000; 
    #10 old_index=5'b00010 ; Q=29'b00010_00_000001_00000011_00000000; 
    #10 old_index=5'b00011 ; Q=29'b00011_00_000001_00000100_00000000;
    #10 old_index=5'b00100 ; Q=29'b00100_00_000001_00000100_00000001; 
    #10 old_index=5'b00101 ; Q=29'b00101_00_000001_00000101_00000100; 
    #10 old_index=5'b00110 ; Q=29'b00110_00_000001_00000110_00000000; 
    #10 old_index=5'b00111 ; Q=29'b00111_00_000001_00000111_00000000;
    #10 old_index=5'b01000 ; Q=29'b01000_00_000001_00001001_00000000; 
    #10 old_index=5'b01001 ; Q=29'b01001_00_000001_00001001_00000111;
    #10 old_index=5'b01010 ; Q=29'b01010_00_000001_00001011_00000000;
    #10 old_index=5'b01011 ; Q=29'b01011_00_000001_00001100_00000000;
    #10 old_index=5'b01100 ; Q=29'b01100_00_000001_00001110_00000000;
    #10 old_index=5'b01101 ; Q=29'b01101_01_000001_00000001_00000000;
    #10 old_index=5'b01110 ; Q=29'b01110_01_000001_00000010_00000000;
    #10 old_index=5'b01111 ; Q=29'b01111_01_000001_00000100_00000000;
    #10 old_index=5'b10000 ; Q=29'b10000_01_000001_00000100_00000001;
    #10 old_index=5'b10001 ; Q=29'b10001_01_000001_00000101_00000100;
    #10 old_index=5'b10010 ; Q=29'b10010_01_000001_00000110_00000000;
    #10 old_index=5'b10011 ; Q=29'b10011_01_000001_00000111_00000000;
    #10 old_index=5'b10100 ; Q=29'b10100_01_000001_00001001_00000000;
    #10 old_index=5'b10101 ; Q=29'b10101_01_000001_00001001_00000111;
    #10 old_index=5'b10110 ; Q=29'b10110_01_000001_00001011_00000000;
    #10 old_index=5'b10111 ; Q=29'b10111_01_000001_00001100_00000000;
    #10 old_index=5'b11000 ; Q=29'b11000_10_000001_00000100_00000001;
    #10 old_index=5'b11001 ; Q=29'b11001_10_000001_00000101_00000100;
    #10 old_index=5'b11010 ; Q=29'b11010_10_000001_00000110_00000000;
    #10 old_index=5'b11011 ; Q=29'b11011_10_000001_00000111_00000000;
    #10 old_index=5'b11100 ; Q=29'b11100_10_000001_00001001_00000000;
    #10 old_index=5'b11101 ; Q=29'b11101_10_000001_00001001_00000111;
    #10 old_index=5'b11110 ; Q=29'b11110_10_000001_00001011_00000000;
    #10 old_index=5'b11111 ; Q=29'b11111_10_000001_00001100_00000000;
    
    #10 $finish;
  end

  initial
  $monitor($time,"'ns| \n %b\n %b\n %b\n %b\n %b\n %b\n %b\n %b\n %b\n %b\n %b\n %b\n %b\n %b\n %b\n %b\n %b\n %b\n %b\n %b\n %b\n %b\n %b\n %b\n %b\n %b\n %b\n %b\n %b\n %b\n %b\n %b",s1, s2, s3, s4, s5, s6, s7, s8, s9, s10, s11, s12, s13, s14, s15, s16, s17, s18, s19, s20, s21, s22, s23, s24, s25, s26, s27, s28, s29, s30, s31, s32);
  //$monitor($time,"'ns| %b \n",  asi);


/*initial begin
//$dumpfile("MCD.vcd");
$dumpfile("MCD_syn.vcd");
$dumpvars;
end         */

endmodule